module cli

pub fn say_hi() {
	println('hello from mymodule!')
}